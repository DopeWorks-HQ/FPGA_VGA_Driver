`timescale 1ns/1ps

module vga_sync(

);

endmodule
